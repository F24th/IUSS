magic
tech scmos
timestamp 1669226985
<< electrodecap >>
rect 21 -100 91 -43
rect -79 -115 91 -100
<< ptransistor >>
rect -77 0 -73 4
rect -22 -8 -17 10
rect -11 -8 -6 10
rect 0 -8 5 10
rect 11 -8 16 10
rect 22 -8 27 10
rect 33 -8 38 10
rect 44 -8 49 10
rect 55 -8 60 10
rect 66 -8 71 10
rect 77 -8 82 10
rect -56 -32 -51 -14
rect -45 -32 -40 -14
rect -22 -32 -17 -14
rect -11 -32 -6 -14
rect 0 -32 5 -14
rect 11 -32 16 -14
rect 22 -32 27 -14
rect 33 -32 38 -14
rect 44 -32 49 -14
rect 55 -32 60 -14
rect 66 -32 71 -14
rect 77 -32 82 -14
<< pdiffusion >>
rect -83 0 -82 4
rect -78 0 -77 4
rect -73 0 -72 4
rect -68 0 -67 4
rect -28 -2 -22 10
rect -28 -8 -27 -2
rect -23 -8 -22 -2
rect -17 4 -16 10
rect -12 4 -11 10
rect -17 -8 -11 4
rect -6 -2 0 10
rect -6 -8 -5 -2
rect -1 -8 0 -2
rect 5 4 6 10
rect 10 4 11 10
rect 5 -8 11 4
rect 16 -2 22 10
rect 16 -8 17 -2
rect 21 -8 22 -2
rect 27 4 28 10
rect 32 4 33 10
rect 27 -8 33 4
rect 38 -2 44 10
rect 38 -8 39 -2
rect 43 -8 44 -2
rect 49 4 50 10
rect 54 4 55 10
rect 49 -8 55 4
rect 60 -2 66 10
rect 60 -8 61 -2
rect 65 -8 66 -2
rect 71 4 72 10
rect 76 4 77 10
rect 71 -8 77 4
rect 82 -2 88 10
rect 82 -8 83 -2
rect 87 -8 88 -2
rect -62 -26 -56 -14
rect -62 -32 -61 -26
rect -57 -32 -56 -26
rect -51 -20 -50 -14
rect -46 -20 -45 -14
rect -51 -32 -45 -20
rect -40 -26 -34 -14
rect -40 -32 -39 -26
rect -35 -32 -34 -26
rect -28 -20 -27 -14
rect -23 -20 -22 -14
rect -28 -32 -22 -20
rect -17 -26 -11 -14
rect -17 -32 -16 -26
rect -12 -32 -11 -26
rect -6 -20 -5 -14
rect -1 -20 0 -14
rect -6 -32 0 -20
rect 5 -26 11 -14
rect 5 -32 6 -26
rect 10 -32 11 -26
rect 16 -20 17 -14
rect 21 -20 22 -14
rect 16 -32 22 -20
rect 27 -26 33 -14
rect 27 -32 28 -26
rect 32 -32 33 -26
rect 38 -20 39 -14
rect 43 -20 44 -14
rect 38 -32 44 -20
rect 49 -26 55 -14
rect 49 -32 50 -26
rect 54 -32 55 -26
rect 60 -20 61 -14
rect 65 -20 66 -14
rect 60 -32 66 -20
rect 71 -26 77 -14
rect 71 -32 72 -26
rect 76 -32 77 -26
rect 82 -20 83 -14
rect 87 -20 88 -14
rect 82 -32 88 -20
<< pdcontact >>
rect -82 0 -78 4
rect -72 0 -68 4
rect -27 -8 -23 -2
rect -16 4 -12 10
rect -5 -8 -1 -2
rect 6 4 10 10
rect 17 -8 21 -2
rect 28 4 32 10
rect 39 -8 43 -2
rect 50 4 54 10
rect 61 -8 65 -2
rect 72 4 76 10
rect 83 -8 87 -2
rect -61 -32 -57 -26
rect -50 -20 -46 -14
rect -39 -32 -35 -26
rect -27 -20 -23 -14
rect -16 -32 -12 -26
rect -5 -20 -1 -14
rect 6 -32 10 -26
rect 17 -20 21 -14
rect 28 -32 32 -26
rect 39 -20 43 -14
rect 50 -32 54 -26
rect 61 -20 65 -14
rect 72 -32 76 -26
rect 83 -20 87 -14
<< nsubstratendiff >>
rect -93 23 107 24
rect -93 19 -87 23
rect 101 19 107 23
rect -93 -36 -92 19
rect -88 18 102 19
rect -88 -36 -87 18
rect -93 -37 -87 -36
rect 101 -36 102 18
rect 106 -36 107 19
rect 101 -37 107 -36
<< nsubstratencontact >>
rect -87 19 101 23
rect -92 -36 -88 19
rect 102 -36 106 19
<< polysilicon >>
rect -22 11 96 16
rect -22 10 -17 11
rect -11 10 -6 11
rect 0 10 5 11
rect 11 10 16 11
rect 22 10 27 11
rect 33 10 38 11
rect 44 10 49 11
rect 55 10 60 11
rect 66 10 71 11
rect 77 10 82 11
rect -77 4 -73 9
rect -77 -3 -73 0
rect -56 -14 -51 -12
rect -45 -14 -40 -12
rect -22 -14 -17 -8
rect -11 -14 -6 -8
rect 0 -14 5 -8
rect 11 -14 16 -8
rect 22 -14 27 -8
rect 33 -14 38 -8
rect 44 -14 49 -8
rect 55 -14 60 -8
rect 66 -14 71 -8
rect 77 -14 82 -8
rect -56 -34 -51 -32
rect -56 -38 -55 -34
rect -45 -35 -40 -32
rect -22 -33 -17 -32
rect -51 -38 -40 -35
rect -19 -34 -17 -33
rect -11 -34 -6 -32
rect 0 -34 5 -32
rect 11 -34 16 -32
rect 22 -34 27 -32
rect 33 -34 38 -32
rect 44 -34 49 -32
rect 55 -34 60 -32
rect 66 -34 71 -32
rect 77 -34 82 -32
rect 91 -34 96 11
rect -19 -37 96 -34
rect -22 -38 96 -37
rect -56 -39 -40 -38
rect 16 -95 96 -38
rect -84 -120 96 -95
<< polycontact >>
rect -77 -7 -73 -3
rect -55 -38 -51 -34
rect -23 -37 -19 -33
<< metal1 >>
rect -92 19 -87 23
rect 101 19 106 23
rect -65 10 -56 19
rect -72 6 -56 10
rect -72 4 -68 6
rect -82 -3 -78 0
rect -82 -7 -77 -3
rect -82 -43 -78 -7
rect -65 -9 -56 6
rect -16 11 94 15
rect -16 10 -12 11
rect 6 10 10 11
rect 28 10 32 11
rect 50 10 54 11
rect 72 10 76 11
rect -27 -9 -23 -8
rect -5 -9 -1 -8
rect 17 -9 21 -8
rect 39 -9 43 -8
rect 61 -9 65 -8
rect 83 -9 87 -8
rect -65 -13 87 -9
rect -50 -14 -46 -13
rect -27 -14 -23 -13
rect -5 -14 -1 -13
rect 17 -14 21 -13
rect 39 -14 43 -13
rect 61 -14 65 -13
rect 83 -14 87 -13
rect -61 -34 -57 -32
rect -39 -33 -35 -32
rect -16 -33 -12 -32
rect 6 -33 10 -32
rect 28 -33 32 -32
rect 50 -33 54 -32
rect 72 -33 76 -32
rect 90 -33 94 11
rect -61 -38 -55 -34
rect -39 -37 -23 -33
rect -16 -37 94 -33
rect -61 -43 -57 -38
rect -39 -43 -35 -37
<< end >>
